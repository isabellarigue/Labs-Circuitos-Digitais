library ieee;
use ieee.std_logic_1164.all;

entity bin2bcd is
	-- Converte um binario (8-bits) para decimal BCD.
	port (
		bin:		in std_logic_vector(7 downto 0);
		dec, un:	out std_logic_vector(3 downto 0)
	);
end;

architecture rtl of bin2bcd is
begin
	-- Utilizacao de tecnicas de programacao orientada a gambiarra (POG)
	with bin select
		un <= "0000" when "00000000",
			"0001" when "00000001",
			"0010" when "00000010",
			"0011" when "00000011",
			"0100" when "00000100",
			"0101" when "00000101",
			"0110" when "00000110",
			"0111" when "00000111",
			"1000" when "00001000",
			"1001" when "00001001",
			"0000" when "00001010",
			"0001" when "00001011",
			"0010" when "00001100",
			"0011" when "00001101",
			"0100" when "00001110",
			"0101" when "00001111",
			"0110" when "00010000",
			"0111" when "00010001",
			"1000" when "00010010",
			"1001" when "00010011",
			"0000" when "00010100",
			"0001" when "00010101",
			"0010" when "00010110",
			"0011" when "00010111",
			"0100" when "00011000",
			"0101" when "00011001",
			"0110" when "00011010",
			"0111" when "00011011",
			"1000" when "00011100",
			"1001" when "00011101",
			"0000" when "00011110",
			"0001" when "00011111",
			"0010" when "00100000",
			"0011" when "00100001",
			"0100" when "00100010",
			"0101" when "00100011",
			"0110" when "00100100",
			"0111" when "00100101",
			"1000" when "00100110",
			"1001" when "00100111",
			"0000" when "00101000",
			"0001" when "00101001",
			"0010" when "00101010",
			"0011" when "00101011",
			"0100" when "00101100",
			"0101" when "00101101",
			"0110" when "00101110",
			"0111" when "00101111",
			"1000" when "00110000",
			"1001" when "00110001",
			"0000" when "00110010",
			"0001" when "00110011",
			"0010" when "00110100",
			"0011" when "00110101",
			"0100" when "00110110",
			"0101" when "00110111",
			"0110" when "00111000",
			"0111" when "00111001",
			"1000" when "00111010",
			"1001" when "00111011",
			"0000" when "00111100",
			"0001" when "00111101",
			"0010" when "00111110",
			"0011" when "00111111",
			"0100" when "01000000",
			"0101" when "01000001",
			"0110" when "01000010",
			"0111" when "01000011",
			"1000" when "01000100",
			"1001" when "01000101",
			"0000" when "01000110",
			"0001" when "01000111",
			"0010" when "01001000",
			"0011" when "01001001",
			"0100" when "01001010",
			"0101" when "01001011",
			"0110" when "01001100",
			"0111" when "01001101",
			"1000" when "01001110",
			"1001" when "01001111",
			"0000" when "01010000",
			"0001" when "01010001",
			"0010" when "01010010",
			"0011" when "01010011",
			"0100" when "01010100",
			"0101" when "01010101",
			"0110" when "01010110",
			"0111" when "01010111",
			"1000" when "01011000",
			"1001" when "01011001",
			"0000" when "01011010",
			"0001" when "01011011",
			"0010" when "01011100",
			"0011" when "01011101",
			"0100" when "01011110",
			"0101" when "01011111",
			"0110" when "01100000",
			"0111" when "01100001",
			"1000" when "01100010",
			"1001" when "01100011",
			"0000" when "01100100",
			"0001" when "01100101",
			"0010" when "01100110",
			"0011" when "01100111",
			"0100" when "01101000",
			"0101" when "01101001",
			"0110" when "01101010",
			"0111" when "01101011",
			"1000" when "01101100",
			"1001" when "01101101",
			"0000" when "01101110",
			"0001" when "01101111",
			"0010" when "01110000",
			"0011" when "01110001",
			"0100" when "01110010",
			"0101" when "01110011",
			"0110" when "01110100",
			"0111" when "01110101",
			"1000" when "01110110",
			"1001" when "01110111",
			"0000" when "01111000",
			"0001" when "01111001",
			"0010" when "01111010",
			"0011" when "01111011",
			"0100" when "01111100",
			"0101" when "01111101",
			"0110" when "01111110",
			"0111" when "01111111",
			"1000" when "10000000",
			"1001" when "10000001",
			"0000" when "10000010",
			"0001" when "10000011",
			"0010" when "10000100",
			"0011" when "10000101",
			"0100" when "10000110",
			"0101" when "10000111",
			"0110" when "10001000",
			"0111" when "10001001",
			"1000" when "10001010",
			"1001" when "10001011",
			"0000" when "10001100",
			"0001" when "10001101",
			"0010" when "10001110",
			"0011" when "10001111",
			"0100" when "10010000",
			"0101" when "10010001",
			"0110" when "10010010",
			"0111" when "10010011",
			"1000" when "10010100",
			"1001" when "10010101",
			"0000" when "10010110",
			"0001" when "10010111",
			"0010" when "10011000",
			"0011" when "10011001",
			"0100" when "10011010",
			"0101" when "10011011",
			"0110" when "10011100",
			"0111" when "10011101",
			"1000" when "10011110",
			"1001" when "10011111",
			"0000" when "10100000",
			"0001" when "10100001",
			"0010" when "10100010",
			"0011" when "10100011",
			"0100" when "10100100",
			"0101" when "10100101",
			"0110" when "10100110",
			"0111" when "10100111",
			"1000" when "10101000",
			"1001" when "10101001",
			"0000" when "10101010",
			"0001" when "10101011",
			"0010" when "10101100",
			"0011" when "10101101",
			"0100" when "10101110",
			"0101" when "10101111",
			"0110" when "10110000",
			"0111" when "10110001",
			"1000" when "10110010",
			"1001" when "10110011",
			"0000" when "10110100",
			"0001" when "10110101",
			"0010" when "10110110",
			"0011" when "10110111",
			"0100" when "10111000",
			"0101" when "10111001",
			"0110" when "10111010",
			"0111" when "10111011",
			"1000" when "10111100",
			"1001" when "10111101",
			"0000" when "10111110",
			"0001" when "10111111",
			"0010" when "11000000",
			"0011" when "11000001",
			"0100" when "11000010",
			"0101" when "11000011",
			"0110" when "11000100",
			"0111" when "11000101",
			"1000" when "11000110",
			"1001" when "11000111",
			"0000" when "11001000",
			"0001" when "11001001",
			"0010" when "11001010",
			"0011" when "11001011",
			"0100" when "11001100",
			"0101" when "11001101",
			"0110" when "11001110",
			"0111" when "11001111",
			"1000" when "11010000",
			"1001" when "11010001",
			"0000" when "11010010",
			"0001" when "11010011",
			"0010" when "11010100",
			"0011" when "11010101",
			"0100" when "11010110",
			"0101" when "11010111",
			"0110" when "11011000",
			"0111" when "11011001",
			"1000" when "11011010",
			"1001" when "11011011",
			"0000" when "11011100",
			"0001" when "11011101",
			"0010" when "11011110",
			"0011" when "11011111",
			"0100" when "11100000",
			"0101" when "11100001",
			"0110" when "11100010",
			"0111" when "11100011",
			"1000" when "11100100",
			"1001" when "11100101",
			"0000" when "11100110",
			"0001" when "11100111",
			"0010" when "11101000",
			"0011" when "11101001",
			"0100" when "11101010",
			"0101" when "11101011",
			"0110" when "11101100",
			"0111" when "11101101",
			"1000" when "11101110",
			"1001" when "11101111",
			"0000" when "11110000",
			"0001" when "11110001",
			"0010" when "11110010",
			"0011" when "11110011",
			"0100" when "11110100",
			"0101" when "11110101",
			"0110" when "11110110",
			"0111" when "11110111",
			"1000" when "11111000",
			"1001" when "11111001",
			"0000" when "11111010",
			"0001" when "11111011",
			"0010" when "11111100",
			"0011" when "11111101",
			"0100" when "11111110",
			"0101" when "11111111",
			"0000" when others;
			
	with bin select
		dec <= "0000" when "00000000",
			"0000" when "00000001",
			"0000" when "00000010",
			"0000" when "00000011",
			"0000" when "00000100",
			"0000" when "00000101",
			"0000" when "00000110",
			"0000" when "00000111",
			"0000" when "00001000",
			"0000" when "00001001",
			"0001" when "00001010",
			"0001" when "00001011",
			"0001" when "00001100",
			"0001" when "00001101",
			"0001" when "00001110",
			"0001" when "00001111",
			"0001" when "00010000",
			"0001" when "00010001",
			"0001" when "00010010",
			"0001" when "00010011",
			"0010" when "00010100",
			"0010" when "00010101",
			"0010" when "00010110",
			"0010" when "00010111",
			"0010" when "00011000",
			"0010" when "00011001",
			"0010" when "00011010",
			"0010" when "00011011",
			"0010" when "00011100",
			"0010" when "00011101",
			"0011" when "00011110",
			"0011" when "00011111",
			"0011" when "00100000",
			"0011" when "00100001",
			"0011" when "00100010",
			"0011" when "00100011",
			"0011" when "00100100",
			"0011" when "00100101",
			"0011" when "00100110",
			"0011" when "00100111",
			"0100" when "00101000",
			"0100" when "00101001",
			"0100" when "00101010",
			"0100" when "00101011",
			"0100" when "00101100",
			"0100" when "00101101",
			"0100" when "00101110",
			"0100" when "00101111",
			"0100" when "00110000",
			"0100" when "00110001",
			"0101" when "00110010",
			"0101" when "00110011",
			"0101" when "00110100",
			"0101" when "00110101",
			"0101" when "00110110",
			"0101" when "00110111",
			"0101" when "00111000",
			"0101" when "00111001",
			"0101" when "00111010",
			"0101" when "00111011",
			"0110" when "00111100",
			"0110" when "00111101",
			"0110" when "00111110",
			"0110" when "00111111",
			"0110" when "01000000",
			"0110" when "01000001",
			"0110" when "01000010",
			"0110" when "01000011",
			"0110" when "01000100",
			"0110" when "01000101",
			"0111" when "01000110",
			"0111" when "01000111",
			"0111" when "01001000",
			"0111" when "01001001",
			"0111" when "01001010",
			"0111" when "01001011",
			"0111" when "01001100",
			"0111" when "01001101",
			"0111" when "01001110",
			"0111" when "01001111",
			"1000" when "01010000",
			"1000" when "01010001",
			"1000" when "01010010",
			"1000" when "01010011",
			"1000" when "01010100",
			"1000" when "01010101",
			"1000" when "01010110",
			"1000" when "01010111",
			"1000" when "01011000",
			"1000" when "01011001",
			"1001" when "01011010",
			"1001" when "01011011",
			"1001" when "01011100",
			"1001" when "01011101",
			"1001" when "01011110",
			"1001" when "01011111",
			"1001" when "01100000",
			"1001" when "01100001",
			"1001" when "01100010",
			"1001" when "01100011",
			"0000" when "01100100",
			"0000" when "01100101",
			"0000" when "01100110",
			"0000" when "01100111",
			"0000" when "01101000",
			"0000" when "01101001",
			"0000" when "01101010",
			"0000" when "01101011",
			"0000" when "01101100",
			"0000" when "01101101",
			"0001" when "01101110",
			"0001" when "01101111",
			"0001" when "01110000",
			"0001" when "01110001",
			"0001" when "01110010",
			"0001" when "01110011",
			"0001" when "01110100",
			"0001" when "01110101",
			"0001" when "01110110",
			"0001" when "01110111",
			"0010" when "01111000",
			"0010" when "01111001",
			"0010" when "01111010",
			"0010" when "01111011",
			"0010" when "01111100",
			"0010" when "01111101",
			"0010" when "01111110",
			"0010" when "01111111",
			"0010" when "10000000",
			"0010" when "10000001",
			"0011" when "10000010",
			"0011" when "10000011",
			"0011" when "10000100",
			"0011" when "10000101",
			"0011" when "10000110",
			"0011" when "10000111",
			"0011" when "10001000",
			"0011" when "10001001",
			"0011" when "10001010",
			"0011" when "10001011",
			"0100" when "10001100",
			"0100" when "10001101",
			"0100" when "10001110",
			"0100" when "10001111",
			"0100" when "10010000",
			"0100" when "10010001",
			"0100" when "10010010",
			"0100" when "10010011",
			"0100" when "10010100",
			"0100" when "10010101",
			"0101" when "10010110",
			"0101" when "10010111",
			"0101" when "10011000",
			"0101" when "10011001",
			"0101" when "10011010",
			"0101" when "10011011",
			"0101" when "10011100",
			"0101" when "10011101",
			"0101" when "10011110",
			"0101" when "10011111",
			"0110" when "10100000",
			"0110" when "10100001",
			"0110" when "10100010",
			"0110" when "10100011",
			"0110" when "10100100",
			"0110" when "10100101",
			"0110" when "10100110",
			"0110" when "10100111",
			"0110" when "10101000",
			"0110" when "10101001",
			"0111" when "10101010",
			"0111" when "10101011",
			"0111" when "10101100",
			"0111" when "10101101",
			"0111" when "10101110",
			"0111" when "10101111",
			"0111" when "10110000",
			"0111" when "10110001",
			"0111" when "10110010",
			"0111" when "10110011",
			"1000" when "10110100",
			"1000" when "10110101",
			"1000" when "10110110",
			"1000" when "10110111",
			"1000" when "10111000",
			"1000" when "10111001",
			"1000" when "10111010",
			"1000" when "10111011",
			"1000" when "10111100",
			"1000" when "10111101",
			"1001" when "10111110",
			"1001" when "10111111",
			"1001" when "11000000",
			"1001" when "11000001",
			"1001" when "11000010",
			"1001" when "11000011",
			"1001" when "11000100",
			"1001" when "11000101",
			"1001" when "11000110",
			"1001" when "11000111",
			"0000" when "11001000",
			"0000" when "11001001",
			"0000" when "11001010",
			"0000" when "11001011",
			"0000" when "11001100",
			"0000" when "11001101",
			"0000" when "11001110",
			"0000" when "11001111",
			"0000" when "11010000",
			"0000" when "11010001",
			"0001" when "11010010",
			"0001" when "11010011",
			"0001" when "11010100",
			"0001" when "11010101",
			"0001" when "11010110",
			"0001" when "11010111",
			"0001" when "11011000",
			"0001" when "11011001",
			"0001" when "11011010",
			"0001" when "11011011",
			"0010" when "11011100",
			"0010" when "11011101",
			"0010" when "11011110",
			"0010" when "11011111",
			"0010" when "11100000",
			"0010" when "11100001",
			"0010" when "11100010",
			"0010" when "11100011",
			"0010" when "11100100",
			"0010" when "11100101",
			"0011" when "11100110",
			"0011" when "11100111",
			"0011" when "11101000",
			"0011" when "11101001",
			"0011" when "11101010",
			"0011" when "11101011",
			"0011" when "11101100",
			"0011" when "11101101",
			"0011" when "11101110",
			"0011" when "11101111",
			"0100" when "11110000",
			"0100" when "11110001",
			"0100" when "11110010",
			"0100" when "11110011",
			"0100" when "11110100",
			"0100" when "11110101",
			"0100" when "11110110",
			"0100" when "11110111",
			"0100" when "11111000",
			"0100" when "11111001",
			"0101" when "11111010",
			"0101" when "11111011",
			"0101" when "11111100",
			"0101" when "11111101",
			"0101" when "11111110",
			"0101" when "11111111",
			"0000" when others;
end rtl;
